`timescale 1ns / 1ps
/**
Alex Knowlton
Single-port synchronous ROM

In Vivado, give name of init file, not relative path. Vivado will handle the relative pathing

parameters:
    depth: number of bits in address
    width: number of bits in output data
    neuron_type: 1 or 0, 1 for fully-connected, 0 for convolutional
    layer_number: layer identifier
    neuron number: neuron identifier
*/

module ROM_neuron #(parameter depth=3, width=8, neuron_type=0, layer_number=1, neuron_number=0) (
    `ifdef VIVADO
    input  logic reset_i,
    `endif
    input  logic clk_i,
    
    /*
    Uncomment when write mode in layers has been resolved
    `ifndef VIVADO
    input logic wen
    input logic [width-1:0] data_i;
    `endif
    */

    input  logic [depth-1:0] addr_i,
    output logic [width-1:0] data_o
    );

    // TODO: Find out if parameters like this negatively impact synthesis
    localparam ascii_offset = 48;
	localparam logic [7:0] neuron_type_p = neuron_type + ascii_offset;
    localparam logic [7:0] layer_number_p = layer_number + ascii_offset;
    localparam logic [7:0] neuron_number_ones_p = (neuron_number % 10) + ascii_offset;
    localparam logic [7:0] neuron_number_tens_p = ((neuron_number / 10) % 10) + ascii_offset;
    localparam logic [7:0] neuron_number_hundreds_p = ((neuron_number / 100) % 10) + ascii_offset;
    

    // odd logic, but it synthesizes to {"n_n_nnn.mem" where "n" is a parameter as defined above}
    localparam logic [87:0] init_file = {neuron_type_p, 8'h5f, layer_number_p, 8'h5f, neuron_number_hundreds_p, neuron_number_tens_p, neuron_number_ones_p, 32'h2e6d656d};
    `ifdef VIVADO
	ROM_inferred #(
        .ADDR_WIDTH(depth),
        .WORD_SIZE(width),
        .MEM_INIT(init_file)
    ) internal_rom (
        .addr_i,
        .data_o,
        .clk_i,
        .reset_i
    );

    `else
    logic wen;
    logic [width-1:0] data_write;
    // TODO: Uncomment when write mode resolved with layers
    // assign data_write = data_i
    
    // remove these two lines when write mode resolved
    assign wen = 1'b0;
    assign data_write = '0;

    generate
        case (neuron_type)
            0: begin
                sram_16_64_freepdk45 ram (
                    .clk0(clk_i),
                    .csb0(1'b0),
                    .web0(wen),
                    .addr0(addr_i),
                    .din0(data_write),
                    .dout0(data_o)
                );
            end
            1: begin
                // larger sram for build, smaller for testing synthesis/apr flow
                `ifdef TESTING
                sram_16_32_freepdk45 ram (
                `else
                sram_16_512_freepdk45 ram (
                `endif
                    .clk0(clk_i),
                    .csb0(1'b0),
                    .web0(wen),
                    .addr0(addr_i),
                    .din0(data_write),
                    .dout0(data_o)
                );
            end
            2: begin
                // larger sram for build, smaller for testing synthesis/apr flow
                `ifdef TESTING
                sram_21_16_freepdk45 ram (
                `else
                sram_21_256_freepdk45 ram (
                `endif
                    .clk0(clk_i),
                    .csb0(1'b0),
                    .web0(wen),
                    .addr0(addr_i),
                    .din0(data_write),
                    .dout0(data_o)
                );
            end
        endcase
    endgenerate
    `endif
    
endmodule