/**
Alex Knowlton
2/28/2023

fully-connected layer
asserts done when first node is done (since all of them work at the same time this is fine)
*/