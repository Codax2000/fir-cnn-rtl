`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 13.11.2018 17:11:05
// Design Name: 
// Module Name: neuron
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created 
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//`define DEBUG
`include "include.v"

module neuron #(parameter layerNo=0,neuronNo=0,numWeight=784,dataWidth=16,sigmoidSize=5,weightIntWidth=1,actType="relu",biasFile="",weightFile="")(
    input           clk,
    input           rst,
    input [dataWidth-1:0]    myinput,
    input           myinputValid,
    input           weightValid,
    input           biasValid,
    input [31:0]    weightValue,
    input [31:0]    biasValue,
    input [31:0]    config_layer_num,
    input [31:0]    config_neuron_num,
    output[dataWidth-1:0]    out,
    output reg      outvalid   
    );
    
    parameter addressWidth = $clog2(numWeight); //clog2(x) = ceiling[log2(x)] -> num of bits I need to count x weights. (x memory slots)
    
    reg         wen;
    wire        ren;
    reg [addressWidth-1:0] w_addr;
    reg [addressWidth:0]   r_addr;     //read address has to reach until numWeight hence width is 1 bit more
    reg [dataWidth-1:0]  w_in;
    wire [dataWidth-1:0] w_out;
    reg [2*dataWidth-1:0]  mul; 
    reg [2*dataWidth-1:0]  sum;
    reg [2*dataWidth-1:0]  bias;
    reg [31:0]    biasReg[0:0];
    reg         weight_valid;
    reg         mult_valid;
    wire        mux_valid;
    reg         sigValid; 
    wire [2*dataWidth:0] comboAdd;
    wire [2*dataWidth:0] BiasAdd;
    reg  [dataWidth-1:0] myinputd;
    reg muxValid_d;
    reg muxValid_f;
    reg addr=0;

   // ------------------------------------------- Loading weight values into the memory -------------------------------------------
    always @(posedge clk)
    begin
        if(rst)                                 // If rst 
        begin
            w_addr <= {addressWidth{1'b1}};     // w_addr<=[11111...1]
                                                // This way, the first time I write sth (look line 76: w_addr <= w_addr + 1)
                                                // it will be writter on w_addr=[0000...0]
            wen <=0;
        end
        else if(weightValid & (config_layer_num==layerNo) & (config_neuron_num==neuronNo))     // when valid weight is comming 
                                                                                               // & layerNo and neuronNo have been defined
        begin
            w_in <= weightValue;        // weight value goes to weight memory
            w_addr <= w_addr + 1;       // all 3 commands happen @ the same time so the weight is written in w_addr + 1
            wen <= 1;
        end
        else
            wen <= 0;
    end

    // --------------------------------------- Dettermine pretrained or not ----------------------------------------
    assign mux_valid = mult_valid;
    assign comboAdd = mul + sum;
    assign BiasAdd = bias + sum;
    assign ren = myinputValid;
    
    `ifdef pretrained
        initial
        begin
            $readmemb(biasFile,biasReg);
        end
        always @(posedge clk)
        begin
            bias <= {biasReg[addr][dataWidth-1:0],{dataWidth{1'b0}}};
        end
    `else
        always @(posedge clk)
        begin
            if(biasValid & (config_layer_num==layerNo) & (config_neuron_num==neuronNo))
            begin
                bias <= {biasValue[dataWidth-1:0],{dataWidth{1'b0}}};
            end
        end
    `endif
    
   // ------------------------------------------- Moving r_addr pointer -------------------------------------------
    always @(posedge clk)
    begin
        if(rst|outvalid)        // -------------- When rst happens OR neuron gives out its output -> raddr is set back to zero ------------
            r_addr <= 0;
        else if(myinputValid)   // NORMAL OPERATION -- Moving to next raddr in next cycle
            r_addr <= r_addr + 1;
    end
    
   // ------------------------------------------- Multiplication -------------------------------------------
    always @(posedge clk)
    begin
        mul  <= $signed(myinputd) * $signed(w_out); // my_input_delayed_by_1_clk * output_of_weight_memory
    end
    
    // -----------------------------------------------------------------------------------------------------
    always @(posedge clk)
    begin
        if(rst|outvalid)        // -------------- When rst happens OR neuron gives out its output -> sum is set back to 0 ------------
            sum <= 0;
        else if((r_addr == numWeight) & muxValid_f) // -------------- if r_addr == max value OR mucValid is falling ----------------
        begin
            if(!bias[2*dataWidth-1] &!sum[2*dataWidth-1] & BiasAdd[2*dataWidth-1]) //If bias and sum are positive and after adding bias to sum, if sign bit becomes 1, saturate
            begin
                sum[2*dataWidth-1] <= 1'b0;
                sum[2*dataWidth-2:0] <= {2*dataWidth-1{1'b1}};
            end
            else if(bias[2*dataWidth-1] & sum[2*dataWidth-1] &  !BiasAdd[2*dataWidth-1]) //If bias and sum are negative and after addition if sign bit is 0, saturate
            begin
                sum[2*dataWidth-1] <= 1'b1;
                sum[2*dataWidth-2:0] <= {2*dataWidth-1{1'b0}};
            end
            else
                sum <= BiasAdd; 
        end
        else if(mux_valid)          // ------------------ NORMAL OPERRATION ------------------
        begin
            if(!mul[2*dataWidth-1] & !sum[2*dataWidth-1] & comboAdd[2*dataWidth-1])  // !mul[2*dataWidth-1] = MSB of mul
                                                                                     // MSB of mul and sum == 0 && MSB of their addition == 1
                                                                                     // meanning we add 2 pos numbers and we get 1 negative
                                                                                     // OVERFLOW
                                                                                     // saturate the output
            begin
                sum[2*dataWidth-1] <= 1'b0;                         // MSB <= 0 (to have a possitive number)
                sum[2*dataWidth-2:0] <= {2*dataWidth-1{1'b1}};      // all rest bits are "1" -> saturation (max num I can get)
            end
            else if(mul[2*dataWidth-1] & sum[2*dataWidth-1] & !comboAdd[2*dataWidth-1])  // UNDERFLOW (neg + neg = pos)
            begin
                sum[2*dataWidth-1] <= 1'b1;                     // MSB <= 1 (to have a negative number)
                sum[2*dataWidth-2:0] <= {2*dataWidth-1{1'b0}};  // all rest bits are "0" -> saturation (min num I can get)
                                                                // remember for -1111 i will write 0_0000 -> the bits are inverted
            end
            else
                sum <= comboAdd; // neither overflow nor underflow
        end
    end
    
   // ------------------------------------------- Loading weight values into the memory ------------------------------------------
    // data is loaded sequentially to each neuron (if I have 5 inputs I neep 5 cucles to read them)
    always @(posedge clk)
    begin
        myinputd <= myinput;                                                // input delayed by 1 clk
        weight_valid <= myinputValid;
        mult_valid <= weight_valid;
        sigValid <= ((r_addr == numWeight) & muxValid_f) ? 1'b1 : 1'b0;
        outvalid <= sigValid;
        muxValid_d <= mux_valid;
        muxValid_f <= !mux_valid & muxValid_d;
    end
        
    // ------------------------------------------- Instantiation of Memory for Weights -------------------------------------------
    Weight_Memory #(.numWeight(numWeight),.neuronNo(neuronNo),.layerNo(layerNo),.addressWidth(addressWidth),.dataWidth(dataWidth),.weightFile(weightFile)) WM(
        .clk(clk),
        .wen(wen),
        .ren(ren),
        .wadd(w_addr),
        .radd(r_addr),
        .win(w_in),
        .wout(w_out)
    );
    
    // ----------------------------- generate statement to selectively instantiate one of the modules -----------------------------------
    generate
        if(actType == "sigmoid")
        begin:siginst
        //Instantiation of ROM for sigmoid
            Sig_ROM #(.inWidth(sigmoidSize),.dataWidth(dataWidth)) s1(
            .clk(clk),
            .x(sum[2*dataWidth-1-:sigmoidSize]),
            .out(out)
        );
        end
        else
        begin:ReLUinst
            ReLU #(.dataWidth(dataWidth),.weightIntWidth(weightIntWidth)) s1 (
            .clk(clk),
            .x(sum),
            .out(out)
        );
        end
    endgenerate

    // ----------------------------- DEBUGGING PRINTS -----------------------------------
    `ifdef DEBUG
    always @(posedge clk)
    begin
        if(outvalid)
            $display(neuronNo,,,,"%b",out);
    end
    `endif

endmodule
