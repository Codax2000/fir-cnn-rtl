module bn_layer_tb ();

endmodule